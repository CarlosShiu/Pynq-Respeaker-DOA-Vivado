`define    AXIS_TDATA_W    32
`define    AXIL_DATA_W     32
`define    AB4C_ADDR_W     12
`define    ENABLE          1
`define    DISABLE         0
`define    RESET_ENABLE_   0